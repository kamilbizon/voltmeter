`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 11/25/2019 01:45:09 PM
// Design Name: 
// Module Name: sterowanie
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


//module sterowanie(
//    input clk,
//    input rst, en,
//    output [7:0] data_rec,
    
//    //ADC side
//    input data1,
//    output cs,
//    output sck
//    );
    
//always @(posedge clk, posedge rst)
//    if(rst)
        
//    else
    
//endmodule
